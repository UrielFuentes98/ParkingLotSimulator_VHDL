LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_BIT.ALL;


ENTITY CLK20HZ IS
	PORT (
		MCLK : IN BIT;
		CLKOUT : OUT BIT);
END CLK20HZ;

ARCHITECTURE Behavioral OF CLK20HZ IS
	SIGNAL COUNTER : INTEGER RANGE 0 TO 250_000 := 0;
	SIGNAL C20HZ: BIT;
BEGIN
	
	PROCESS (MCLK)
	BEGIN
		IF MCLK = '1' AND MCLK'EVENT THEN
			IF COUNTER = 250_000 THEN
				COUNTER <= 0;
				C20HZ <= NOT C20HZ;
			ELSE COUNTER <= COUNTER + 1;
		END IF;
		ELSE NULL;
		END IF;
	END PROCESS;
				 CLKOUT <= C20HZ ;
				 
END Behavioral;